----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:27:03 11/06/2018 
-- Design Name: 
-- Module Name:    SSegDisplay - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
--                        a
--                      =====
--                    b|| g ||f
--                      =====
--                    c||   ||e
--                      =====
--                        d  
-- ____________________________________________________________________
-- |iCNT0|iCNT1|iCNT2|iCNT3||  a  |  b  |  c  |  d  |  e  |  f  |  g  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  0  |  0  |  0  |  0  ||  1  |  1  |  1  |  1  |  1  |  1  |  0  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  0  |  0  |  0  |  1  ||  0  |  0  |  0  |  0  |  1  |  1  |  0  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  0  |  0  |  1  |  0  ||  1  |  0  |  1  |  1  |  0  |  1  |  1  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  0  |  0  |  1  |  1  ||  1  |  1  |  0  |  0  |  1  |  1  |  1  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  0  |  1  |  0  |  0  ||  0  |  1  |  0  |  0  |  1  |  1  |  1  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  0  |  1  |  0  |  1  ||  1  |  1  |  0  |  1  |  1  |  0  |  1  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  0  |  1  |  1  |  0  ||  1  |  1  |  1  |  1  |  1  |  0  |  1  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  0  |  1  |  1  |  1  ||  1  |  0  |  0  |  0  |  1  |  1  |  0  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  1  |  0  |  0  |  0  ||  1  |  1  |  1  |  1  |  1  |  1  |  1  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  1  |  0  |  0  |  1  ||  1  |  1  |  0  |  1  |  1  |  1  |  1  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  1  |  0  |  1  |  0  ||  1  |  1  |  1  |  0  |  1  |  1  |  1  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  1  |  0  |  1  |  1  ||  0  |  1  |  1  |  1  |  1  |  0  |  1  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  1  |  1  |  0  |  0  ||  1  |  1  |  1  |  1  |  0  |  0  |  0  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  1  |  1  |  0  |  1  ||  0  |  0  |  1  |  1  |  1  |  1  |  1  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  1  |  1  |  1  |  0  ||  1  |  1  |  1  |  1  |  0  |  0  |  1  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
-- |  1  |  1  |  1  |  1  ||  1  |  1  |  1  |  0  |  0  |  0  |  1  |
-- |_____|_____|_____|_____||_____|_____|_____|_____|_____|_____|_____|
--
-- oSSeg(6:0) = (a, b, c, d, e, f, g)   

-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SSegDisplay is
    Port ( iCNT  : in  std_logic_vector(3 downto 0);
           oSSeg : out std_logic_vector(6 downto 0));
end SSegDisplay;

architecture Behavioral of SSegDisplay is
     
begin
    with iCNT select oSSeg <=
	     "1111110" when "0000",
	     "0000110" when "0001",
	     "1111010" when "0010",
	     "1100110" when "0011",
	     "0100101" when "0100",
	     "1101101" when "0101",
	     "1011111" when "0110",
	     "1100110" when "0111",
	     "1111111" when "1000",
	     "1101111" when "1001",
	     "1110111" when "1010",
	     "0111101" when "1011",
	     "1111000" when "1100",
	     "0011111" when "1101",
	     "1111001" when "1110",
	     "1110001" when "1111",
	     "0110111" when others;		  

end Behavioral;

